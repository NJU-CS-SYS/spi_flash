module SPIFlashModule(input clk, input reset,
    input  io_flash_en,
    input  io_flash_write,
    input [3:0] io_quad_io,
    input [23:0] io_flash_addr,
    input [31:0] io_flash_data_in,
    output[31:0] io_flash_data_out,
    output[11:0] io_state_to_cpu,
    output io_SI,
    output io_tri_si,
    output io_cs,
    output io_ready
);

  reg  cs;
  wire T401;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire not_move;
  wire T11;
  wire T12;
  reg  write_old;
  wire T402;
  wire T13;
  wire T14;
  reg [5:0] state;
  wire[5:0] T403;
  wire[5:0] T15;
  wire[5:0] T16;
  wire[5:0] T17;
  wire[5:0] T18;
  wire[5:0] T19;
  wire[5:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg [5:0] counter;
  wire[5:0] T404;
  wire[6:0] T405;
  wire[6:0] T32;
  wire[6:0] T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  wire[6:0] T406;
  wire[5:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire[5:0] T46;
  wire[5:0] T47;
  wire[5:0] T48;
  wire[5:0] T49;
  wire[5:0] T50;
  wire[5:0] T51;
  wire[5:0] T52;
  wire[5:0] T53;
  wire[5:0] T54;
  wire[5:0] T55;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire[5:0] T59;
  wire[5:0] T60;
  wire[5:0] T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire[5:0] T65;
  wire[5:0] T66;
  wire[5:0] T67;
  wire[5:0] T68;
  wire[5:0] T69;
  wire T70;
  wire T71;
  reg [5:0] sub_state;
  wire[5:0] T407;
  wire[5:0] T72;
  wire[5:0] T73;
  wire[5:0] T74;
  wire[5:0] T75;
  wire[5:0] T76;
  wire[5:0] T77;
  wire[5:0] T78;
  wire[5:0] T79;
  wire[5:0] T80;
  wire[5:0] T81;
  wire[5:0] T82;
  wire[5:0] T83;
  wire[5:0] T84;
  wire[5:0] T85;
  wire[5:0] T86;
  wire[5:0] T87;
  wire[5:0] T88;
  wire[5:0] T89;
  wire[5:0] T90;
  wire[5:0] T91;
  wire[5:0] T92;
  wire[5:0] T93;
  wire[5:0] T94;
  wire[5:0] T95;
  wire[5:0] T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire[5:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[5:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[5:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire[5:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[5:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire[5:0] T131;
  wire T132;
  wire T133;
  wire[5:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[5:0] T139;
  wire[5:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire[5:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire[5:0] T151;
  wire T152;
  wire T153;
  wire[5:0] T154;
  wire T155;
  wire T156;
  wire[5:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[5:0] T162;
  wire T163;
  wire T164;
  wire[5:0] T165;
  wire[5:0] T166;
  wire[5:0] T408;
  wire[3:0] T167;
  wire[3:0] T168;
  wire[1:0] T409;
  wire T410;
  wire[5:0] T169;
  wire[5:0] T170;
  wire[5:0] T171;
  wire[5:0] T172;
  wire[6:0] T173;
  wire[6:0] T174;
  wire[6:0] T175;
  wire[6:0] T411;
  wire T176;
  wire T177;
  wire[6:0] T178;
  wire[6:0] T179;
  wire[6:0] T412;
  wire T180;
  wire T181;
  wire[6:0] T182;
  wire[6:0] T413;
  wire[2:0] T183;
  wire[2:0] T184;
  wire[2:0] T185;
  wire[2:0] T186;
  wire[6:0] T187;
  wire[6:0] T414;
  wire[3:0] T188;
  wire[3:0] T189;
  wire[2:0] T415;
  wire T416;
  wire T190;
  wire T191;
  wire[6:0] T192;
  wire[6:0] T417;
  wire[4:0] T193;
  wire[1:0] T194;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[6:0] T197;
  wire[6:0] T418;
  wire[5:0] T198;
  wire[5:0] T199;
  wire T419;
  wire T200;
  wire T201;
  wire[2:0] T202;
  wire[6:0] T420;
  wire[5:0] T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  reg [23:0] addr_old;
  wire[23:0] T421;
  wire[23:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[1:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire[2:0] T262;
  reg [7:0] RDCR;
  wire[7:0] T422;
  wire T263;
  wire[2:0] T264;
  reg [7:0] RDSR1;
  wire[7:0] T423;
  wire T265;
  wire[2:0] T266;
  reg [7:0] WRR;
  wire[7:0] T424;
  wire T267;
  wire[2:0] T268;
  reg [7:0] reg_buffer_sr1;
  wire[7:0] T425;
  wire[8:0] T426;
  wire[8:0] T269;
  wire[8:0] T270;
  wire[8:0] T427;
  wire[8:0] T271;
  wire[8:0] T272;
  wire[8:0] T273;
  wire[8:0] T274;
  wire[7:0] T275;
  wire[2:0] T276;
  wire[8:0] T428;
  wire T277;
  wire T278;
  wire T279;
  wire[8:0] T280;
  wire[8:0] T281;
  wire[8:0] T429;
  wire[8:0] T282;
  wire[8:0] T283;
  wire[8:0] T284;
  wire[8:0] T285;
  wire[7:0] T286;
  wire[2:0] T287;
  wire[8:0] T430;
  wire T288;
  wire T289;
  wire T290;
  wire[8:0] T291;
  wire[8:0] T292;
  wire T293;
  wire[2:0] T294;
  reg [7:0] reg_buffer_cr;
  wire[7:0] T431;
  wire[8:0] T432;
  wire[8:0] T295;
  wire[8:0] T296;
  wire[8:0] T433;
  wire[8:0] T297;
  wire[8:0] T298;
  wire[8:0] T299;
  wire[8:0] T300;
  wire[7:0] T301;
  wire[2:0] T302;
  wire[8:0] T434;
  wire T303;
  wire T304;
  wire T305;
  wire[8:0] T306;
  wire[8:0] T307;
  wire[8:0] T435;
  wire[8:0] T436;
  wire[7:0] T308;
  wire T309;
  wire[2:0] T310;
  wire T311;
  wire[2:0] T312;
  reg [7:0] QREAD;
  wire[7:0] T437;
  wire T313;
  wire[4:0] T314;
  wire T315;
  wire[2:0] T316;
  reg [7:0] WREN;
  wire[7:0] T438;
  wire T317;
  wire[2:0] T318;
  reg [7:0] PP;
  wire[7:0] T439;
  wire T319;
  wire[4:0] T320;
  wire T321;
  wire[4:0] T322;
  wire T323;
  wire[2:0] T324;
  wire[11:0] T325;
  reg [31:0] buffer;
  wire[31:0] T440;
  wire[32:0] T441;
  wire[32:0] T326;
  wire[32:0] T327;
  wire[32:0] T442;
  wire[31:0] T328;
  wire[31:0] T329;
  wire[31:0] T330;
  wire[31:0] T331;
  wire[31:0] T332;
  wire[31:0] T333;
  wire[31:0] T334;
  wire[31:0] T443;
  wire[7:0] T335;
  wire[3:0] T336;
  wire[31:0] T337;
  wire[31:0] T444;
  wire[8:0] T338;
  wire[8:0] T339;
  wire[22:0] T445;
  wire T446;
  wire T340;
  wire[31:0] T341;
  wire[31:0] T447;
  wire[3:0] T342;
  wire[3:0] T343;
  wire[31:0] T344;
  wire[31:0] T448;
  wire[4:0] T345;
  wire[4:0] T346;
  wire[26:0] T449;
  wire T450;
  wire T347;
  wire T348;
  wire T349;
  wire[31:0] T350;
  wire[31:0] T451;
  wire[15:0] T351;
  wire[3:0] T352;
  wire[31:0] T353;
  wire[31:0] T452;
  wire[16:0] T354;
  wire[16:0] T355;
  wire[14:0] T453;
  wire T454;
  wire T356;
  wire T357;
  wire T358;
  wire[31:0] T359;
  wire[31:0] T455;
  wire[11:0] T360;
  wire[3:0] T361;
  wire[31:0] T362;
  wire[31:0] T456;
  wire[12:0] T363;
  wire[12:0] T364;
  wire[18:0] T457;
  wire T458;
  wire T365;
  wire T366;
  wire T367;
  wire[31:0] T368;
  wire[31:0] T459;
  wire[23:0] T369;
  wire[3:0] T370;
  wire[31:0] T371;
  wire[31:0] T460;
  wire[24:0] T372;
  wire[24:0] T373;
  wire[6:0] T461;
  wire T462;
  wire T374;
  wire T375;
  wire T376;
  wire[31:0] T377;
  wire[31:0] T463;
  wire[19:0] T378;
  wire[3:0] T379;
  wire[31:0] T380;
  wire[31:0] T464;
  wire[20:0] T381;
  wire[20:0] T382;
  wire[10:0] T465;
  wire T466;
  wire T383;
  wire T384;
  wire T385;
  wire[32:0] T386;
  wire[32:0] T467;
  wire[31:0] T387;
  wire[3:0] T388;
  wire[32:0] T389;
  wire[32:0] T390;
  wire[32:0] T391;
  wire[32:0] T468;
  wire T392;
  wire T393;
  wire T394;
  wire[32:0] T395;
  wire[32:0] T469;
  wire[27:0] T396;
  wire[3:0] T397;
  wire[32:0] T398;
  wire[32:0] T470;
  wire[28:0] T399;
  wire[28:0] T400;
  wire[3:0] T471;
  wire T472;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    cs = {1{$random}};
    write_old = {1{$random}};
    state = {1{$random}};
    counter = {1{$random}};
    sub_state = {1{$random}};
    addr_old = {1{$random}};
    RDCR = {1{$random}};
    RDSR1 = {1{$random}};
    WRR = {1{$random}};
    reg_buffer_sr1 = {1{$random}};
    reg_buffer_cr = {1{$random}};
    QREAD = {1{$random}};
    WREN = {1{$random}};
    PP = {1{$random}};
    buffer = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_ready = {1{$random}};
// synthesis translate_on
`endif
  assign io_cs = cs;
  assign T401 = reset ? 1'h1 : T0;
  assign T0 = T245 ? 1'h1 : T1;
  assign T1 = T243 ? 1'h0 : T2;
  assign T2 = T241 ? 1'h1 : T3;
  assign T3 = T226 ? 1'h1 : T4;
  assign T4 = T224 ? 1'h0 : T5;
  assign T5 = T222 ? 1'h1 : T6;
  assign T6 = T220 ? 1'h0 : T7;
  assign T7 = T218 ? 1'h0 : T8;
  assign T8 = T9 ? 1'h0 : cs;
  assign T9 = T217 & T10;
  assign T10 = ~ not_move;
  assign not_move = T214 | T11;
  assign T11 = T210 & T12;
  assign T12 = write_old == io_flash_write;
  assign T402 = reset ? 1'h0 : T13;
  assign T13 = T14 ? io_flash_write : write_old;
  assign T14 = state == 6'h3;
  assign T403 = reset ? 6'h0 : T15;
  assign T15 = T14 ? 6'h0 : T16;
  assign T16 = T245 ? 6'h3 : T17;
  assign T17 = T226 ? 6'h3 : T18;
  assign T18 = T26 ? 6'h1 : T19;
  assign T19 = T24 ? 6'h2 : T20;
  assign T20 = T21 ? 6'h4 : state;
  assign T21 = T9 & T22;
  assign T22 = io_flash_en & T23;
  assign T23 = ~ io_flash_write;
  assign T24 = T9 & T25;
  assign T25 = io_flash_en & io_flash_write;
  assign T26 = T30 & T27;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T29 == 1'h1;
  assign T29 = io_quad_io[1];
  assign T30 = T208 & T31;
  assign T31 = counter == 6'h0;
  assign T404 = T405[5:0];
  assign T405 = reset ? 7'h0 : T32;
  assign T32 = T206 ? 7'h7 : T33;
  assign T33 = T204 ? T420 : T34;
  assign T34 = T245 ? 7'h7 : T35;
  assign T35 = T200 ? T192 : T36;
  assign T36 = T190 ? T182 : T37;
  assign T37 = T180 ? T173 : T406;
  assign T406 = {1'h0, T38};
  assign T38 = T180 ? T169 : T39;
  assign T39 = T180 ? T165 : T40;
  assign T40 = T163 ? T162 : T41;
  assign T41 = T160 ? 6'h17 : T42;
  assign T42 = T158 ? T157 : T43;
  assign T43 = T241 ? 6'h7 : T44;
  assign T44 = T155 ? T154 : T45;
  assign T45 = T152 ? T151 : T46;
  assign T46 = T149 ? 6'h0 : T47;
  assign T47 = T147 ? T146 : T48;
  assign T48 = T144 ? 6'h17 : T49;
  assign T49 = T141 ? T140 : T50;
  assign T50 = T26 ? 6'h7 : T51;
  assign T51 = T208 ? T139 : T52;
  assign T52 = T137 ? 6'h7 : T53;
  assign T53 = T135 ? T134 : T54;
  assign T54 = T222 ? 6'h7 : T55;
  assign T55 = T132 ? T131 : T56;
  assign T56 = T129 ? 6'h7 : T57;
  assign T57 = T127 ? T126 : T58;
  assign T58 = T124 ? 6'h7 : T59;
  assign T59 = T122 ? T121 : T60;
  assign T60 = T119 ? 6'h7 : T61;
  assign T61 = T117 ? T116 : T62;
  assign T62 = T114 ? 6'h7 : T63;
  assign T63 = T112 ? T111 : T64;
  assign T64 = T109 ? 6'h7 : T65;
  assign T65 = T107 ? T106 : T66;
  assign T66 = T104 ? 6'h7 : T67;
  assign T67 = T70 ? T69 : T68;
  assign T68 = T9 ? 6'h7 : counter;
  assign T69 = counter - 6'h1;
  assign T70 = T103 & T71;
  assign T71 = sub_state == 6'hb;
  assign T407 = reset ? 6'h0 : T72;
  assign T72 = T98 ? 6'h9 : T73;
  assign T73 = T206 ? 6'ha : T74;
  assign T74 = T245 ? 6'h0 : T75;
  assign T75 = T180 ? 6'h8 : T76;
  assign T76 = T160 ? 6'h5 : T77;
  assign T77 = T243 ? 6'h4 : T78;
  assign T78 = T241 ? 6'h7 : T79;
  assign T79 = T226 ? 6'h0 : T80;
  assign T80 = T149 ? 6'h6 : T81;
  assign T81 = T144 ? 6'h5 : T82;
  assign T82 = T26 ? 6'h4 : T83;
  assign T83 = T97 ? 6'h10 : T84;
  assign T84 = T137 ? 6'h11 : T85;
  assign T85 = T224 ? 6'h10 : T86;
  assign T86 = T222 ? 6'h13 : T87;
  assign T87 = T129 ? 6'hf : T88;
  assign T88 = T124 ? 6'he : T89;
  assign T89 = T220 ? 6'hd : T90;
  assign T90 = T119 ? 6'h12 : T91;
  assign T91 = T114 ? 6'ha : T92;
  assign T92 = T218 ? 6'h3 : T93;
  assign T93 = T109 ? 6'h7 : T94;
  assign T94 = T104 ? 6'hc : T95;
  assign T95 = T24 ? 6'h1 : T96;
  assign T96 = T21 ? 6'hb : sub_state;
  assign T97 = T30 & T28;
  assign T98 = T100 & T99;
  assign T99 = counter == 6'h0;
  assign T100 = T102 & T101;
  assign T101 = sub_state == 6'ha;
  assign T102 = state == 6'h2;
  assign T103 = state == 6'h4;
  assign T104 = T70 & T105;
  assign T105 = counter == 6'h0;
  assign T106 = counter - 6'h1;
  assign T107 = T103 & T108;
  assign T108 = sub_state == 6'hc;
  assign T109 = T107 & T110;
  assign T110 = counter == 6'h0;
  assign T111 = counter - 6'h1;
  assign T112 = T103 & T113;
  assign T113 = sub_state == 6'h3;
  assign T114 = T112 & T115;
  assign T115 = counter == 6'h0;
  assign T116 = counter - 6'h1;
  assign T117 = T103 & T118;
  assign T118 = sub_state == 6'ha;
  assign T119 = T117 & T120;
  assign T120 = counter == 6'h0;
  assign T121 = counter - 6'h1;
  assign T122 = T103 & T123;
  assign T123 = sub_state == 6'hd;
  assign T124 = T122 & T125;
  assign T125 = counter == 6'h0;
  assign T126 = counter - 6'h1;
  assign T127 = T103 & T128;
  assign T128 = sub_state == 6'he;
  assign T129 = T127 & T130;
  assign T130 = counter == 6'h0;
  assign T131 = counter - 6'h1;
  assign T132 = T103 & T133;
  assign T133 = sub_state == 6'hf;
  assign T134 = counter - 6'h1;
  assign T135 = T103 & T136;
  assign T136 = sub_state == 6'h10;
  assign T137 = T135 & T138;
  assign T138 = counter == 6'h0;
  assign T139 = counter - 6'h1;
  assign T140 = counter - 6'h1;
  assign T141 = T143 & T142;
  assign T142 = sub_state == 6'h4;
  assign T143 = state == 6'h1;
  assign T144 = T141 & T145;
  assign T145 = counter == 6'h0;
  assign T146 = counter - 6'h1;
  assign T147 = T143 & T148;
  assign T148 = sub_state == 6'h5;
  assign T149 = T147 & T150;
  assign T150 = counter == 6'h0;
  assign T151 = counter + 6'h1;
  assign T152 = T143 & T153;
  assign T153 = sub_state == 6'h6;
  assign T154 = counter - 6'h1;
  assign T155 = T102 & T156;
  assign T156 = sub_state == 6'h1;
  assign T157 = counter - 6'h1;
  assign T158 = T102 & T159;
  assign T159 = sub_state == 6'h4;
  assign T160 = T158 & T161;
  assign T161 = counter == 6'h0;
  assign T162 = counter - 6'h1;
  assign T163 = T102 & T164;
  assign T164 = sub_state == 6'h5;
  assign T165 = T166 | 6'h7;
  assign T166 = T40 & T408;
  assign T408 = {T409, T167};
  assign T167 = ~ T168;
  assign T168 = 4'h7;
  assign T409 = T410 ? 2'h3 : 2'h0;
  assign T410 = T167[3];
  assign T169 = T170 | 6'h0;
  assign T170 = T39 & T171;
  assign T171 = ~ T172;
  assign T172 = 6'h18;
  assign T173 = T178 | T174;
  assign T174 = T411 & T175;
  assign T175 = 7'h20;
  assign T411 = T176 ? 7'h7f : 7'h0;
  assign T176 = T177;
  assign T177 = 1'h0;
  assign T178 = T412 & T179;
  assign T179 = ~ T175;
  assign T412 = {1'h0, T38};
  assign T180 = T163 & T181;
  assign T181 = counter == 6'h0;
  assign T182 = T187 | T413;
  assign T413 = {4'h0, T183};
  assign T183 = T184 << 1'h0;
  assign T184 = T185 & 3'h7;
  assign T185 = T186 - 3'h1;
  assign T186 = counter[2:0];
  assign T187 = T37 & T414;
  assign T414 = {T415, T188};
  assign T188 = ~ T189;
  assign T189 = 4'h7;
  assign T415 = T416 ? 3'h7 : 3'h0;
  assign T416 = T188[3];
  assign T190 = T102 & T191;
  assign T191 = sub_state == 6'h8;
  assign T192 = T197 | T417;
  assign T417 = {2'h0, T193};
  assign T193 = T194 << 2'h3;
  assign T194 = T195 & 2'h3;
  assign T195 = T196 + 2'h1;
  assign T196 = counter[4:3];
  assign T197 = T36 & T418;
  assign T418 = {T419, T198};
  assign T198 = ~ T199;
  assign T199 = 6'h18;
  assign T419 = T198[5];
  assign T200 = T190 & T201;
  assign T201 = T202 == 3'h0;
  assign T202 = counter[2:0];
  assign T420 = {1'h0, T203};
  assign T203 = counter - 6'h1;
  assign T204 = T102 & T205;
  assign T205 = sub_state == 6'h3;
  assign T206 = T204 & T207;
  assign T207 = counter == 6'h0;
  assign T208 = T103 & T209;
  assign T209 = sub_state == 6'h11;
  assign T210 = T213 & T211;
  assign T211 = addr_old == io_flash_addr;
  assign T421 = reset ? 24'h0 : T212;
  assign T212 = T14 ? io_flash_addr : addr_old;
  assign T213 = state == 6'h0;
  assign T214 = T216 & T215;
  assign T215 = io_flash_en == 1'h0;
  assign T216 = state == 6'h0;
  assign T217 = state == 6'h0;
  assign T218 = T103 & T219;
  assign T219 = sub_state == 6'h7;
  assign T220 = T103 & T221;
  assign T221 = sub_state == 6'h12;
  assign T222 = T132 & T223;
  assign T223 = counter == 6'h0;
  assign T224 = T103 & T225;
  assign T225 = sub_state == 6'h13;
  assign T226 = T152 & T227;
  assign T227 = T228 ^ 1'h1;
  assign T228 = T230 | T229;
  assign T229 = counter == 6'h6;
  assign T230 = T232 | T231;
  assign T231 = counter == 6'h5;
  assign T232 = T234 | T233;
  assign T233 = counter == 6'h4;
  assign T234 = T236 | T235;
  assign T235 = counter == 6'h3;
  assign T236 = T238 | T237;
  assign T237 = counter == 6'h2;
  assign T238 = T240 | T239;
  assign T239 = counter == 6'h1;
  assign T240 = counter == 6'h0;
  assign T241 = T155 & T242;
  assign T242 = counter == 6'h0;
  assign T243 = T102 & T244;
  assign T244 = sub_state == 6'h7;
  assign T245 = T200 & T246;
  assign T246 = T247 == 2'h3;
  assign T247 = counter[4:3];
  assign io_tri_si = T152;
  assign io_SI = T248;
  assign T248 = T204 ? T323 : T249;
  assign T249 = T190 ? T321 : T250;
  assign T250 = T163 ? T319 : T251;
  assign T251 = T158 ? T317 : T252;
  assign T252 = T155 ? T315 : T253;
  assign T253 = T147 ? T313 : T254;
  assign T254 = T141 ? T311 : T255;
  assign T255 = T135 ? T309 : T256;
  assign T256 = T132 ? T293 : T257;
  assign T257 = T127 ? T267 : T258;
  assign T258 = T122 ? T265 : T259;
  assign T259 = T112 ? T263 : T260;
  assign T260 = T70 ? T261 : 1'h0;
  assign T261 = RDCR[T262];
  assign T262 = counter[2:0];
  assign T422 = reset ? 8'h35 : RDCR;
  assign T263 = RDSR1[T264];
  assign T264 = counter[2:0];
  assign T423 = reset ? 8'h5 : RDSR1;
  assign T265 = WRR[T266];
  assign T266 = counter[2:0];
  assign T424 = reset ? 8'h1 : WRR;
  assign T267 = reg_buffer_sr1[T268];
  assign T268 = counter[2:0];
  assign T425 = T426[7:0];
  assign T426 = reset ? 9'h0 : T269;
  assign T269 = T208 ? T282 : T270;
  assign T270 = T117 ? T271 : T427;
  assign T427 = {1'h0, reg_buffer_sr1};
  assign T271 = T280 | T272;
  assign T272 = T428 & T273;
  assign T273 = T274;
  assign T274 = {1'h0, T275};
  assign T275 = 1'h1 << T276;
  assign T276 = counter[2:0];
  assign T428 = T277 ? 9'h1ff : 9'h0;
  assign T277 = T278;
  assign T278 = T279;
  assign T279 = io_quad_io[1];
  assign T280 = T429 & T281;
  assign T281 = ~ T273;
  assign T429 = {1'h0, reg_buffer_sr1};
  assign T282 = T291 | T283;
  assign T283 = T430 & T284;
  assign T284 = T285;
  assign T285 = {1'h0, T286};
  assign T286 = 1'h1 << T287;
  assign T287 = counter[2:0];
  assign T430 = T288 ? 9'h1ff : 9'h0;
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = io_quad_io[1];
  assign T291 = T270 & T292;
  assign T292 = ~ T284;
  assign T293 = reg_buffer_cr[T294];
  assign T294 = counter[2:0];
  assign T431 = T432[7:0];
  assign T432 = reset ? 9'h0 : T295;
  assign T295 = T129 ? T436 : T296;
  assign T296 = T107 ? T297 : T433;
  assign T433 = {1'h0, reg_buffer_cr};
  assign T297 = T306 | T298;
  assign T298 = T434 & T299;
  assign T299 = T300;
  assign T300 = {1'h0, T301};
  assign T301 = 1'h1 << T302;
  assign T302 = counter[2:0];
  assign T434 = T303 ? 9'h1ff : 9'h0;
  assign T303 = T304;
  assign T304 = T305;
  assign T305 = io_quad_io[1];
  assign T306 = T435 & T307;
  assign T307 = ~ T299;
  assign T435 = {1'h0, reg_buffer_cr};
  assign T436 = {1'h0, T308};
  assign T308 = reg_buffer_cr | 8'h2;
  assign T309 = RDSR1[T310];
  assign T310 = counter[2:0];
  assign T311 = QREAD[T312];
  assign T312 = counter[2:0];
  assign T437 = reset ? 8'h6b : QREAD;
  assign T313 = io_flash_addr[T314];
  assign T314 = counter[4:0];
  assign T315 = WREN[T316];
  assign T316 = counter[2:0];
  assign T438 = reset ? 8'h6 : WREN;
  assign T317 = PP[T318];
  assign T318 = counter[2:0];
  assign T439 = reset ? 8'h2 : PP;
  assign T319 = io_flash_addr[T320];
  assign T320 = counter[4:0];
  assign T321 = io_flash_data_in[T322];
  assign T322 = counter[4:0];
  assign T323 = RDSR1[T324];
  assign T324 = counter[2:0];
  assign io_state_to_cpu = T325;
  assign T325 = {state, sub_state};
  assign io_flash_data_out = buffer;
  assign T440 = T441[31:0];
  assign T441 = reset ? 33'h0 : T326;
  assign T326 = T226 ? T395 : T327;
  assign T327 = T392 ? T386 : T442;
  assign T442 = {1'h0, T328};
  assign T328 = T383 ? T377 : T329;
  assign T329 = T374 ? T368 : T330;
  assign T330 = T365 ? T359 : T331;
  assign T331 = T356 ? T350 : T332;
  assign T332 = T347 ? T341 : T333;
  assign T333 = T340 ? T334 : buffer;
  assign T334 = T337 | T443;
  assign T443 = {24'h0, T335};
  assign T335 = T336 << 3'h4;
  assign T336 = io_quad_io & 4'hf;
  assign T337 = buffer & T444;
  assign T444 = {T445, T338};
  assign T338 = ~ T339;
  assign T339 = 9'hf0;
  assign T445 = T446 ? 23'h7fffff : 23'h0;
  assign T446 = T338[8];
  assign T340 = T152 & T240;
  assign T341 = T344 | T447;
  assign T447 = {28'h0, T342};
  assign T342 = T343 << 1'h0;
  assign T343 = io_quad_io & 4'hf;
  assign T344 = T333 & T448;
  assign T448 = {T449, T345};
  assign T345 = ~ T346;
  assign T346 = 5'hf;
  assign T449 = T450 ? 27'h7ffffff : 27'h0;
  assign T450 = T345[4];
  assign T347 = T152 & T348;
  assign T348 = T349 & T239;
  assign T349 = T240 ^ 1'h1;
  assign T350 = T353 | T451;
  assign T451 = {16'h0, T351};
  assign T351 = T352 << 4'hc;
  assign T352 = io_quad_io & 4'hf;
  assign T353 = T332 & T452;
  assign T452 = {T453, T354};
  assign T354 = ~ T355;
  assign T355 = 17'hf000;
  assign T453 = T454 ? 15'h7fff : 15'h0;
  assign T454 = T354[16];
  assign T356 = T152 & T357;
  assign T357 = T358 & T237;
  assign T358 = T238 ^ 1'h1;
  assign T359 = T362 | T455;
  assign T455 = {20'h0, T360};
  assign T360 = T361 << 4'h8;
  assign T361 = io_quad_io & 4'hf;
  assign T362 = T331 & T456;
  assign T456 = {T457, T363};
  assign T363 = ~ T364;
  assign T364 = 13'hf00;
  assign T457 = T458 ? 19'h7ffff : 19'h0;
  assign T458 = T363[12];
  assign T365 = T152 & T366;
  assign T366 = T367 & T235;
  assign T367 = T236 ^ 1'h1;
  assign T368 = T371 | T459;
  assign T459 = {8'h0, T369};
  assign T369 = T370 << 5'h14;
  assign T370 = io_quad_io & 4'hf;
  assign T371 = T330 & T460;
  assign T460 = {T461, T372};
  assign T372 = ~ T373;
  assign T373 = 25'hf00000;
  assign T461 = T462 ? 7'h7f : 7'h0;
  assign T462 = T372[24];
  assign T374 = T152 & T375;
  assign T375 = T376 & T233;
  assign T376 = T234 ^ 1'h1;
  assign T377 = T380 | T463;
  assign T463 = {12'h0, T378};
  assign T378 = T379 << 5'h10;
  assign T379 = io_quad_io & 4'hf;
  assign T380 = T329 & T464;
  assign T464 = {T465, T381};
  assign T381 = ~ T382;
  assign T382 = 21'hf0000;
  assign T465 = T466 ? 11'h7ff : 11'h0;
  assign T466 = T381[20];
  assign T383 = T152 & T384;
  assign T384 = T385 & T231;
  assign T385 = T232 ^ 1'h1;
  assign T386 = T389 | T467;
  assign T467 = {1'h0, T387};
  assign T387 = T388 << 5'h1c;
  assign T388 = io_quad_io & 4'hf;
  assign T389 = T468 & T390;
  assign T390 = ~ T391;
  assign T391 = 33'hf0000000;
  assign T468 = {1'h0, T328};
  assign T392 = T152 & T393;
  assign T393 = T394 & T229;
  assign T394 = T230 ^ 1'h1;
  assign T395 = T398 | T469;
  assign T469 = {5'h0, T396};
  assign T396 = T397 << 5'h18;
  assign T397 = io_quad_io & 4'hf;
  assign T398 = T327 & T470;
  assign T470 = {T471, T399};
  assign T399 = ~ T400;
  assign T400 = 29'hf000000;
  assign T471 = T472 ? 4'hf : 4'h0;
  assign T472 = T399[28];

  always @(posedge clk) begin
    if(reset) begin
      cs <= 1'h1;
    end else if(T245) begin
      cs <= 1'h1;
    end else if(T243) begin
      cs <= 1'h0;
    end else if(T241) begin
      cs <= 1'h1;
    end else if(T226) begin
      cs <= 1'h1;
    end else if(T224) begin
      cs <= 1'h0;
    end else if(T222) begin
      cs <= 1'h1;
    end else if(T220) begin
      cs <= 1'h0;
    end else if(T218) begin
      cs <= 1'h0;
    end else if(T9) begin
      cs <= 1'h0;
    end
    if(reset) begin
      write_old <= 1'h0;
    end else if(T14) begin
      write_old <= io_flash_write;
    end
    if(reset) begin
      state <= 6'h0;
    end else if(T14) begin
      state <= 6'h0;
    end else if(T245) begin
      state <= 6'h3;
    end else if(T226) begin
      state <= 6'h3;
    end else if(T26) begin
      state <= 6'h1;
    end else if(T24) begin
      state <= 6'h2;
    end else if(T21) begin
      state <= 6'h4;
    end
    counter <= T404;
    if(reset) begin
      sub_state <= 6'h0;
    end else if(T98) begin
      sub_state <= 6'h9;
    end else if(T206) begin
      sub_state <= 6'ha;
    end else if(T245) begin
      sub_state <= 6'h0;
    end else if(T180) begin
      sub_state <= 6'h8;
    end else if(T160) begin
      sub_state <= 6'h5;
    end else if(T243) begin
      sub_state <= 6'h4;
    end else if(T241) begin
      sub_state <= 6'h7;
    end else if(T226) begin
      sub_state <= 6'h0;
    end else if(T149) begin
      sub_state <= 6'h6;
    end else if(T144) begin
      sub_state <= 6'h5;
    end else if(T26) begin
      sub_state <= 6'h4;
    end else if(T97) begin
      sub_state <= 6'h10;
    end else if(T137) begin
      sub_state <= 6'h11;
    end else if(T224) begin
      sub_state <= 6'h10;
    end else if(T222) begin
      sub_state <= 6'h13;
    end else if(T129) begin
      sub_state <= 6'hf;
    end else if(T124) begin
      sub_state <= 6'he;
    end else if(T220) begin
      sub_state <= 6'hd;
    end else if(T119) begin
      sub_state <= 6'h12;
    end else if(T114) begin
      sub_state <= 6'ha;
    end else if(T218) begin
      sub_state <= 6'h3;
    end else if(T109) begin
      sub_state <= 6'h7;
    end else if(T104) begin
      sub_state <= 6'hc;
    end else if(T24) begin
      sub_state <= 6'h1;
    end else if(T21) begin
      sub_state <= 6'hb;
    end
    if(reset) begin
      addr_old <= 24'h0;
    end else if(T14) begin
      addr_old <= io_flash_addr;
    end
    if(reset) begin
      RDCR <= 8'h35;
    end
    if(reset) begin
      RDSR1 <= 8'h5;
    end
    if(reset) begin
      WRR <= 8'h1;
    end
    reg_buffer_sr1 <= T425;
    reg_buffer_cr <= T431;
    if(reset) begin
      QREAD <= 8'h6b;
    end
    if(reset) begin
      WREN <= 8'h6;
    end
    if(reset) begin
      PP <= 8'h2;
    end
    buffer <= T440;
  end
endmodule

