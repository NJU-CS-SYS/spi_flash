module SPIFlashModule(input clk, input reset,
    input  io_flash_en,
    input  io_flash_write,
    input [3:0] io_quad_io,
    input [23:0] io_flash_addr,
    input [31:0] io_flash_data_in,
    output[31:0] io_flash_data_out,
    output[11:0] io_state_to_cpu,
    output io_SI,
    output io_tri_si,
    output io_cs
);

  reg  cs;
  wire T252;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire not_move;
  wire T7;
  wire T8;
  reg  write_old;
  wire T253;
  wire T9;
  wire T10;
  reg [5:0] state;
  wire[5:0] T254;
  wire[5:0] T11;
  wire[5:0] T12;
  wire[5:0] T13;
  wire[5:0] T14;
  wire[5:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  reg [23:0] addr_old;
  wire[23:0] T255;
  wire[23:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg [5:0] counter;
  wire[5:0] T256;
  wire[6:0] T257;
  wire[6:0] T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T258;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire[5:0] T46;
  wire[5:0] T47;
  wire[5:0] T48;
  wire[5:0] T49;
  wire[5:0] T50;
  wire[5:0] T51;
  wire[5:0] T52;
  wire T53;
  wire T54;
  reg [5:0] sub_state;
  wire[5:0] T259;
  wire[5:0] T55;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire[5:0] T59;
  wire[5:0] T60;
  wire[5:0] T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire[5:0] T65;
  wire[5:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[5:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[5:0] T80;
  wire[5:0] T81;
  wire T82;
  wire T83;
  wire[5:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire[5:0] T89;
  wire T90;
  wire T91;
  wire[5:0] T92;
  wire[5:0] T93;
  wire[5:0] T260;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[1:0] T261;
  wire T262;
  wire[5:0] T96;
  wire[5:0] T97;
  wire[5:0] T98;
  wire[5:0] T99;
  wire[6:0] T100;
  wire[6:0] T101;
  wire[6:0] T102;
  wire[6:0] T263;
  wire T103;
  wire T104;
  wire[6:0] T105;
  wire[6:0] T106;
  wire[6:0] T264;
  wire T107;
  wire T108;
  wire[6:0] T109;
  wire[6:0] T265;
  wire[2:0] T110;
  wire[2:0] T111;
  wire[2:0] T112;
  wire[2:0] T113;
  wire[6:0] T114;
  wire[6:0] T266;
  wire[3:0] T115;
  wire[3:0] T116;
  wire[2:0] T267;
  wire T268;
  wire T117;
  wire T118;
  wire[6:0] T119;
  wire[6:0] T269;
  wire[4:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[6:0] T124;
  wire[6:0] T270;
  wire[5:0] T125;
  wire[5:0] T126;
  wire T271;
  wire T127;
  wire T128;
  wire[2:0] T129;
  wire[6:0] T272;
  wire[5:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire[1:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[2:0] T163;
  reg [7:0] QREAD;
  wire[7:0] T273;
  wire T164;
  wire[4:0] T165;
  wire T166;
  wire[2:0] T167;
  reg [7:0] WREN;
  wire[7:0] T274;
  wire T168;
  wire[2:0] T169;
  reg [7:0] PP;
  wire[7:0] T275;
  wire T170;
  wire[4:0] T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire[2:0] T175;
  reg [7:0] RDSR1;
  wire[7:0] T276;
  wire[11:0] T176;
  reg [31:0] buffer;
  wire[31:0] T277;
  wire[32:0] T278;
  wire[32:0] T177;
  wire[32:0] T178;
  wire[32:0] T279;
  wire[31:0] T179;
  wire[31:0] T180;
  wire[31:0] T181;
  wire[31:0] T182;
  wire[31:0] T183;
  wire[31:0] T184;
  wire[31:0] T185;
  wire[31:0] T280;
  wire[7:0] T186;
  wire[3:0] T187;
  wire[31:0] T188;
  wire[31:0] T281;
  wire[8:0] T189;
  wire[8:0] T190;
  wire[22:0] T282;
  wire T283;
  wire T191;
  wire[31:0] T192;
  wire[31:0] T284;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[31:0] T195;
  wire[31:0] T285;
  wire[4:0] T196;
  wire[4:0] T197;
  wire[26:0] T286;
  wire T287;
  wire T198;
  wire T199;
  wire T200;
  wire[31:0] T201;
  wire[31:0] T288;
  wire[15:0] T202;
  wire[3:0] T203;
  wire[31:0] T204;
  wire[31:0] T289;
  wire[16:0] T205;
  wire[16:0] T206;
  wire[14:0] T290;
  wire T291;
  wire T207;
  wire T208;
  wire T209;
  wire[31:0] T210;
  wire[31:0] T292;
  wire[11:0] T211;
  wire[3:0] T212;
  wire[31:0] T213;
  wire[31:0] T293;
  wire[12:0] T214;
  wire[12:0] T215;
  wire[18:0] T294;
  wire T295;
  wire T216;
  wire T217;
  wire T218;
  wire[31:0] T219;
  wire[31:0] T296;
  wire[23:0] T220;
  wire[3:0] T221;
  wire[31:0] T222;
  wire[31:0] T297;
  wire[24:0] T223;
  wire[24:0] T224;
  wire[6:0] T298;
  wire T299;
  wire T225;
  wire T226;
  wire T227;
  wire[31:0] T228;
  wire[31:0] T300;
  wire[19:0] T229;
  wire[3:0] T230;
  wire[31:0] T231;
  wire[31:0] T301;
  wire[20:0] T232;
  wire[20:0] T233;
  wire[10:0] T302;
  wire T303;
  wire T234;
  wire T235;
  wire T236;
  wire[32:0] T237;
  wire[32:0] T304;
  wire[31:0] T238;
  wire[3:0] T239;
  wire[32:0] T240;
  wire[32:0] T241;
  wire[32:0] T242;
  wire[32:0] T305;
  wire T243;
  wire T244;
  wire T245;
  wire[32:0] T246;
  wire[32:0] T306;
  wire[27:0] T247;
  wire[3:0] T248;
  wire[32:0] T249;
  wire[32:0] T307;
  wire[28:0] T250;
  wire[28:0] T251;
  wire[3:0] T308;
  wire T309;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    cs = {1{$random}};
    write_old = {1{$random}};
    state = {1{$random}};
    addr_old = {1{$random}};
    counter = {1{$random}};
    sub_state = {1{$random}};
    QREAD = {1{$random}};
    WREN = {1{$random}};
    PP = {1{$random}};
    RDSR1 = {1{$random}};
    buffer = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_cs = cs;
  assign T252 = reset ? 1'h1 : T0;
  assign T0 = T152 ? 1'h1 : T1;
  assign T1 = T150 ? 1'h0 : T2;
  assign T2 = T148 ? 1'h1 : T3;
  assign T3 = T29 ? 1'h1 : T4;
  assign T4 = T5 ? 1'h0 : cs;
  assign T5 = T28 & T6;
  assign T6 = ~ not_move;
  assign not_move = T25 | T7;
  assign T7 = T21 & T8;
  assign T8 = write_old == io_flash_write;
  assign T253 = reset ? 1'h0 : T9;
  assign T9 = T10 ? io_flash_write : write_old;
  assign T10 = state == 6'h3;
  assign T254 = reset ? 6'h0 : T11;
  assign T11 = T10 ? 6'h0 : T12;
  assign T12 = T152 ? 6'h3 : T13;
  assign T13 = T29 ? 6'h3 : T14;
  assign T14 = T19 ? 6'h2 : T15;
  assign T15 = T16 ? 6'h1 : state;
  assign T16 = T5 & T17;
  assign T17 = io_flash_en & T18;
  assign T18 = ~ io_flash_write;
  assign T19 = T5 & T20;
  assign T20 = io_flash_en & io_flash_write;
  assign T21 = T24 & T22;
  assign T22 = addr_old == io_flash_addr;
  assign T255 = reset ? 24'h0 : T23;
  assign T23 = T10 ? io_flash_addr : addr_old;
  assign T24 = state == 6'h0;
  assign T25 = T27 & T26;
  assign T26 = io_flash_en == 1'h0;
  assign T27 = state == 6'h0;
  assign T28 = state == 6'h0;
  assign T29 = T146 & T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T135 | T32;
  assign T32 = counter == 6'h6;
  assign T256 = T257[5:0];
  assign T257 = reset ? 7'h0 : T33;
  assign T33 = T133 ? 7'h7 : T34;
  assign T34 = T131 ? T272 : T35;
  assign T35 = T152 ? 7'h7 : T36;
  assign T36 = T127 ? T119 : T37;
  assign T37 = T117 ? T109 : T38;
  assign T38 = T107 ? T100 : T258;
  assign T258 = {1'h0, T39};
  assign T39 = T107 ? T96 : T40;
  assign T40 = T107 ? T92 : T41;
  assign T41 = T90 ? T89 : T42;
  assign T42 = T87 ? 6'h17 : T43;
  assign T43 = T85 ? T84 : T44;
  assign T44 = T148 ? 6'h7 : T45;
  assign T45 = T82 ? T81 : T46;
  assign T46 = T146 ? T80 : T47;
  assign T47 = T78 ? 6'h0 : T48;
  assign T48 = T76 ? T75 : T49;
  assign T49 = T73 ? 6'h17 : T50;
  assign T50 = T53 ? T52 : T51;
  assign T51 = T5 ? 6'h7 : counter;
  assign T52 = counter - 6'h1;
  assign T53 = T72 & T54;
  assign T54 = sub_state == 6'h4;
  assign T259 = reset ? 6'h0 : T55;
  assign T55 = T67 ? 6'h9 : T56;
  assign T56 = T133 ? 6'ha : T57;
  assign T57 = T152 ? 6'h0 : T58;
  assign T58 = T107 ? 6'h8 : T59;
  assign T59 = T87 ? 6'h5 : T60;
  assign T60 = T150 ? 6'h4 : T61;
  assign T61 = T148 ? 6'h7 : T62;
  assign T62 = T29 ? 6'h0 : T63;
  assign T63 = T78 ? 6'h6 : T64;
  assign T64 = T73 ? 6'h5 : T65;
  assign T65 = T19 ? 6'h1 : T66;
  assign T66 = T16 ? 6'h4 : sub_state;
  assign T67 = T69 & T68;
  assign T68 = counter == 6'h0;
  assign T69 = T71 & T70;
  assign T70 = sub_state == 6'ha;
  assign T71 = state == 6'h2;
  assign T72 = state == 6'h1;
  assign T73 = T53 & T74;
  assign T74 = counter == 6'h0;
  assign T75 = counter - 6'h1;
  assign T76 = T72 & T77;
  assign T77 = sub_state == 6'h5;
  assign T78 = T76 & T79;
  assign T79 = counter == 6'h0;
  assign T80 = counter + 6'h1;
  assign T81 = counter - 6'h1;
  assign T82 = T71 & T83;
  assign T83 = sub_state == 6'h1;
  assign T84 = counter - 6'h1;
  assign T85 = T71 & T86;
  assign T86 = sub_state == 6'h4;
  assign T87 = T85 & T88;
  assign T88 = counter == 6'h0;
  assign T89 = counter - 6'h1;
  assign T90 = T71 & T91;
  assign T91 = sub_state == 6'h5;
  assign T92 = T93 | 6'h7;
  assign T93 = T41 & T260;
  assign T260 = {T261, T94};
  assign T94 = ~ T95;
  assign T95 = 4'h7;
  assign T261 = T262 ? 2'h3 : 2'h0;
  assign T262 = T94[3];
  assign T96 = T97 | 6'h0;
  assign T97 = T40 & T98;
  assign T98 = ~ T99;
  assign T99 = 6'h18;
  assign T100 = T105 | T101;
  assign T101 = T263 & T102;
  assign T102 = 7'h20;
  assign T263 = T103 ? 7'h7f : 7'h0;
  assign T103 = T104;
  assign T104 = 1'h0;
  assign T105 = T264 & T106;
  assign T106 = ~ T102;
  assign T264 = {1'h0, T39};
  assign T107 = T90 & T108;
  assign T108 = counter == 6'h0;
  assign T109 = T114 | T265;
  assign T265 = {4'h0, T110};
  assign T110 = T111 << 1'h0;
  assign T111 = T112 & 3'h7;
  assign T112 = T113 - 3'h1;
  assign T113 = counter[2:0];
  assign T114 = T38 & T266;
  assign T266 = {T267, T115};
  assign T115 = ~ T116;
  assign T116 = 4'h7;
  assign T267 = T268 ? 3'h7 : 3'h0;
  assign T268 = T115[3];
  assign T117 = T71 & T118;
  assign T118 = sub_state == 6'h8;
  assign T119 = T124 | T269;
  assign T269 = {2'h0, T120};
  assign T120 = T121 << 2'h3;
  assign T121 = T122 & 2'h3;
  assign T122 = T123 + 2'h1;
  assign T123 = counter[4:3];
  assign T124 = T37 & T270;
  assign T270 = {T271, T125};
  assign T125 = ~ T126;
  assign T126 = 6'h18;
  assign T271 = T125[5];
  assign T127 = T117 & T128;
  assign T128 = T129 == 3'h0;
  assign T129 = counter[2:0];
  assign T272 = {1'h0, T130};
  assign T130 = counter - 6'h1;
  assign T131 = T71 & T132;
  assign T132 = sub_state == 6'h3;
  assign T133 = T131 & T134;
  assign T134 = counter == 6'h0;
  assign T135 = T137 | T136;
  assign T136 = counter == 6'h5;
  assign T137 = T139 | T138;
  assign T138 = counter == 6'h4;
  assign T139 = T141 | T140;
  assign T140 = counter == 6'h3;
  assign T141 = T143 | T142;
  assign T142 = counter == 6'h2;
  assign T143 = T145 | T144;
  assign T144 = counter == 6'h1;
  assign T145 = counter == 6'h0;
  assign T146 = T72 & T147;
  assign T147 = sub_state == 6'h6;
  assign T148 = T82 & T149;
  assign T149 = counter == 6'h0;
  assign T150 = T71 & T151;
  assign T151 = sub_state == 6'h7;
  assign T152 = T127 & T153;
  assign T153 = T154 == 2'h3;
  assign T154 = counter[4:3];
  assign io_tri_si = T146;
  assign io_SI = T155;
  assign T155 = T131 ? T174 : T156;
  assign T156 = T117 ? T172 : T157;
  assign T157 = T90 ? T170 : T158;
  assign T158 = T85 ? T168 : T159;
  assign T159 = T82 ? T166 : T160;
  assign T160 = T76 ? T164 : T161;
  assign T161 = T53 ? T162 : 1'h0;
  assign T162 = QREAD[T163];
  assign T163 = counter[2:0];
  assign T273 = reset ? 8'h6b : QREAD;
  assign T164 = io_flash_addr[T165];
  assign T165 = counter[4:0];
  assign T166 = WREN[T167];
  assign T167 = counter[2:0];
  assign T274 = reset ? 8'h6 : WREN;
  assign T168 = PP[T169];
  assign T169 = counter[2:0];
  assign T275 = reset ? 8'h2 : PP;
  assign T170 = io_flash_addr[T171];
  assign T171 = counter[4:0];
  assign T172 = io_flash_data_in[T173];
  assign T173 = counter[4:0];
  assign T174 = RDSR1[T175];
  assign T175 = counter[2:0];
  assign T276 = reset ? 8'h5 : RDSR1;
  assign io_state_to_cpu = T176;
  assign T176 = {state, sub_state};
  assign io_flash_data_out = buffer;
  assign T277 = T278[31:0];
  assign T278 = reset ? 33'h0 : T177;
  assign T177 = T29 ? T246 : T178;
  assign T178 = T243 ? T237 : T279;
  assign T279 = {1'h0, T179};
  assign T179 = T234 ? T228 : T180;
  assign T180 = T225 ? T219 : T181;
  assign T181 = T216 ? T210 : T182;
  assign T182 = T207 ? T201 : T183;
  assign T183 = T198 ? T192 : T184;
  assign T184 = T191 ? T185 : buffer;
  assign T185 = T188 | T280;
  assign T280 = {24'h0, T186};
  assign T186 = T187 << 3'h4;
  assign T187 = io_quad_io & 4'hf;
  assign T188 = buffer & T281;
  assign T281 = {T282, T189};
  assign T189 = ~ T190;
  assign T190 = 9'hf0;
  assign T282 = T283 ? 23'h7fffff : 23'h0;
  assign T283 = T189[8];
  assign T191 = T146 & T145;
  assign T192 = T195 | T284;
  assign T284 = {28'h0, T193};
  assign T193 = T194 << 1'h0;
  assign T194 = io_quad_io & 4'hf;
  assign T195 = T184 & T285;
  assign T285 = {T286, T196};
  assign T196 = ~ T197;
  assign T197 = 5'hf;
  assign T286 = T287 ? 27'h7ffffff : 27'h0;
  assign T287 = T196[4];
  assign T198 = T146 & T199;
  assign T199 = T200 & T144;
  assign T200 = T145 ^ 1'h1;
  assign T201 = T204 | T288;
  assign T288 = {16'h0, T202};
  assign T202 = T203 << 4'hc;
  assign T203 = io_quad_io & 4'hf;
  assign T204 = T183 & T289;
  assign T289 = {T290, T205};
  assign T205 = ~ T206;
  assign T206 = 17'hf000;
  assign T290 = T291 ? 15'h7fff : 15'h0;
  assign T291 = T205[16];
  assign T207 = T146 & T208;
  assign T208 = T209 & T142;
  assign T209 = T143 ^ 1'h1;
  assign T210 = T213 | T292;
  assign T292 = {20'h0, T211};
  assign T211 = T212 << 4'h8;
  assign T212 = io_quad_io & 4'hf;
  assign T213 = T182 & T293;
  assign T293 = {T294, T214};
  assign T214 = ~ T215;
  assign T215 = 13'hf00;
  assign T294 = T295 ? 19'h7ffff : 19'h0;
  assign T295 = T214[12];
  assign T216 = T146 & T217;
  assign T217 = T218 & T140;
  assign T218 = T141 ^ 1'h1;
  assign T219 = T222 | T296;
  assign T296 = {8'h0, T220};
  assign T220 = T221 << 5'h14;
  assign T221 = io_quad_io & 4'hf;
  assign T222 = T181 & T297;
  assign T297 = {T298, T223};
  assign T223 = ~ T224;
  assign T224 = 25'hf00000;
  assign T298 = T299 ? 7'h7f : 7'h0;
  assign T299 = T223[24];
  assign T225 = T146 & T226;
  assign T226 = T227 & T138;
  assign T227 = T139 ^ 1'h1;
  assign T228 = T231 | T300;
  assign T300 = {12'h0, T229};
  assign T229 = T230 << 5'h10;
  assign T230 = io_quad_io & 4'hf;
  assign T231 = T180 & T301;
  assign T301 = {T302, T232};
  assign T232 = ~ T233;
  assign T233 = 21'hf0000;
  assign T302 = T303 ? 11'h7ff : 11'h0;
  assign T303 = T232[20];
  assign T234 = T146 & T235;
  assign T235 = T236 & T136;
  assign T236 = T137 ^ 1'h1;
  assign T237 = T240 | T304;
  assign T304 = {1'h0, T238};
  assign T238 = T239 << 5'h1c;
  assign T239 = io_quad_io & 4'hf;
  assign T240 = T305 & T241;
  assign T241 = ~ T242;
  assign T242 = 33'hf0000000;
  assign T305 = {1'h0, T179};
  assign T243 = T146 & T244;
  assign T244 = T245 & T32;
  assign T245 = T135 ^ 1'h1;
  assign T246 = T249 | T306;
  assign T306 = {5'h0, T247};
  assign T247 = T248 << 5'h18;
  assign T248 = io_quad_io & 4'hf;
  assign T249 = T178 & T307;
  assign T307 = {T308, T250};
  assign T250 = ~ T251;
  assign T251 = 29'hf000000;
  assign T308 = T309 ? 4'hf : 4'h0;
  assign T309 = T250[28];

  always @(posedge clk) begin
    if(reset) begin
      cs <= 1'h1;
    end else if(T152) begin
      cs <= 1'h1;
    end else if(T150) begin
      cs <= 1'h0;
    end else if(T148) begin
      cs <= 1'h1;
    end else if(T29) begin
      cs <= 1'h1;
    end else if(T5) begin
      cs <= 1'h0;
    end
    if(reset) begin
      write_old <= 1'h0;
    end else if(T10) begin
      write_old <= io_flash_write;
    end
    if(reset) begin
      state <= 6'h0;
    end else if(T10) begin
      state <= 6'h0;
    end else if(T152) begin
      state <= 6'h3;
    end else if(T29) begin
      state <= 6'h3;
    end else if(T19) begin
      state <= 6'h2;
    end else if(T16) begin
      state <= 6'h1;
    end
    if(reset) begin
      addr_old <= 24'h0;
    end else if(T10) begin
      addr_old <= io_flash_addr;
    end
    counter <= T256;
    if(reset) begin
      sub_state <= 6'h0;
    end else if(T67) begin
      sub_state <= 6'h9;
    end else if(T133) begin
      sub_state <= 6'ha;
    end else if(T152) begin
      sub_state <= 6'h0;
    end else if(T107) begin
      sub_state <= 6'h8;
    end else if(T87) begin
      sub_state <= 6'h5;
    end else if(T150) begin
      sub_state <= 6'h4;
    end else if(T148) begin
      sub_state <= 6'h7;
    end else if(T29) begin
      sub_state <= 6'h0;
    end else if(T78) begin
      sub_state <= 6'h6;
    end else if(T73) begin
      sub_state <= 6'h5;
    end else if(T19) begin
      sub_state <= 6'h1;
    end else if(T16) begin
      sub_state <= 6'h4;
    end
    if(reset) begin
      QREAD <= 8'h6b;
    end
    if(reset) begin
      WREN <= 8'h6;
    end
    if(reset) begin
      PP <= 8'h2;
    end
    if(reset) begin
      RDSR1 <= 8'h5;
    end
    buffer <= T277;
  end
endmodule

